module Encoder (
    input clk,
    input rst,
    input [7:0] in_data,
    input in_valid,
    output reg [11:0] out_data,
    output reg out_valid
);



endmodule