module lab7_2(
    input clk,
    input rst,
    input up,
    input down,
    input left,
    input right,
    input hint,
    output [3:0] vgaRed,
    output [3:0] vgaGreen,
    output [3:0] vgaBlue,
    output hsync,
    output vsync,
    output pass
    );
    // add your design here
    
endmodule