`timescale 1ns/100ps
module lab1_2 (
    input wire [5:0] source_0,
    input wire [5:0] source_1,
    input wire [5:0] source_2,
    input wire [5:0] source_3,
    output reg [3:0] result
); 
    /* Note that result can be either reg or wire. 
    * It depends on how you design your module. */
    // add your design here 
endmodule
