module lab3_2
(
    input clk,
    input rst,
    input en,
    input speed,
    input freeze,
    output [15:0] led
);

endmodule
