module Decoder (
    input clk,
    input rst,
    input [11:0] one_bit_err_in_data,
    input one_bit_err_in_valid,
    output reg [7:0] out_plaintext,
    output reg out_plaintext_valid
);



endmodule