module lab3_1
(
    input clk,
    input rst,
    input en,
    input speed,
    output [15:0] led
);

endmodule
