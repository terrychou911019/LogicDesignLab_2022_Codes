module lab7_1(
    input clk,
    input rst,
    input en,
    input dir,
    input vmir,
    input hmir,
    output [3:0] vgaRed,
    output [3:0] vgaGreen,
    output [3:0] vgaBlue,
    output hsync,
    output vsync
);
    // add your design here
    
endmodule